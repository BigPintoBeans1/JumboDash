aoskjd;fkjna;sdf